library verilog;
use verilog.vl_types.all;
entity clk_div_tb is
end clk_div_tb;
