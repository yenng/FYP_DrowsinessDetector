library verilog;
use verilog.vl_types.all;
entity WeightInitialise_tb is
end WeightInitialise_tb;
