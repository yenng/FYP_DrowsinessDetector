module multiply(
input	[9:0] in1,
input	[9:0] in2,
output reg signed [19:0]mulVal
);
reg [9:0] in2_abs,mulVal_t;
//in2 is the value of weight, the data might be negative.

assign mulVal = in1*in2;

//the final answer will be negative if the value of weight is negative. 
//assign mulVal = in2[9] ? -mulVal_t : mulVal_t;
/*module multiply(
input	[9:0] in1,
input	[9:0] in2,
output reg signed [19:0]mulVal
);
reg [9:0] in2_abs,mulVal_t;
//in2 is the value of weight, the data might be negative.
assign in2 = in2 - 10'b1000000000;

//the final answer will be negative if the value of weight is negative. 
assign mulVal = in1*in2;
endmodule*/

endmodule