library verilog;
use verilog.vl_types.all;
entity WeightRAM_sv_unit is
end WeightRAM_sv_unit;
