library verilog;
use verilog.vl_types.all;
entity HiddenLayer_tb is
end HiddenLayer_tb;
