module WeighInitiallize(
	input Clock, In, WE,
	input [3:0] weightNew,
	input [3:0] address,
	output reg weight [0:9][0:9]
);
integer i, seed;
reg [31:0] rand;


endmodule

 