module counter(
	input clk,start,
	input [9:0]max,
	output reg stop,
	output reg[9:0]count
);


always@(posedge clk) begin
	if (start) begin
		if(count == max-1)begin
			stop = 1;
		end
		else begin
			count++;
		end
	end
	else begin
		count = 10'b0;
		stop = 0;
	end
end

endmodule