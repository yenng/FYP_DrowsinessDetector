library verilog;
use verilog.vl_types.all;
entity WeightOptimization_tb is
end WeightOptimization_tb;
