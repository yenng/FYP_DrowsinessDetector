library verilog;
use verilog.vl_types.all;
entity SigmoidPrime_tb is
end SigmoidPrime_tb;
