module HiddenLayer();
	
endmodule 