library verilog;
use verilog.vl_types.all;
entity WeightRAM_tb is
end WeightRAM_tb;
