library verilog;
use verilog.vl_types.all;
entity WeightUpdate_tb is
end WeightUpdate_tb;
