module DrowsinessDetector(
	input Clock,Rst,Start,training,
	input [9:0] in1 [29:0],
	input [9:0] out_ann_real[2:0],
	output reg [9:0] out_ann[2:0],
	output reg [9:0] out_hid[4:0],
	output reg [3:0] state,
	output [9:0]delta1[2:0],
	output [2:0]sign1);
	
	//reg training; // Used to make decision whether train or detect.
	
	// For RAM to write/read weight. 
	reg WE;
	reg signed[9:0]dataOut;
	reg signed[9:0] dataIn;
	
	// The random data that generated by LFSR.
	reg signed[9:0] data;
	reg on;
	
	// The address of RAM to call the weight.
	reg [7:0] Address;
	
	// The variable that represent the state and nextState.
	reg [3:0] nextState;
	
	// Parameter for the state.
	parameter 	halt = 0, weightInitiallize = 1, readWeight = 2, halt1 = 3, hiddenLayer = 4,
	           outputLayer = 5, readWeight1 = 6, halt2 = 7, weightOptimize = 8, weightUpdate = 9,
	           halt0 = 10, writeWeight = 11;
	
	// The variable for hidden layer.
	reg Clear;
	reg signed[9:0]sum;
	reg [9:0]AF_in;
	reg [9:0] AF;
	reg signed [9:0] weight;
	reg unsigned[9:0]inVal;
	reg unsigned[9:0]inVal1;
	reg [9:0] count0,count1;
	reg [9:0] out0[4:0];
	reg [9:0] out1[2:0];
	
	// The variable for weight optimization
	wire [9:0]out1_err[2:0];
	wire [9:0]sig_prime_1[2:0];
	//wire [9:0]delta1[0:2];
	//wire [2:0]sign1;
	
	always@(posedge Clock, negedge Rst) begin
		if(~Rst) begin
			state <= halt0;
		end
		else begin
			state <= nextState;
		end
	end
	
	always@( Start, state, training, data, dataOut) begin
		case(state)
		  // The following state is for weightInitiallize module.
		  halt0: begin 
		    on = 0;
		    Clear = 1;
		    count0 = 0;
		    count1 = 0;
				out0[0] = 10'd0;
				out0[1] = 10'd0;
				out0[2] = 10'd0;
				out0[3] = 10'd0;
				out0[4] = 10'd0;
				out1[0] = 10'd0;
				out1[1] = 10'd0;
				out1[2] = 10'd0;
		    nextState = weightInitiallize;
		  end
			halt: begin
			  WE = 0;
				on = 0;				// Off LFSR
				Address = count0+count1*10'd30;
				if(Start)
					nextState = readWeight;
				else 
				  nextState = halt;
			end
			weightInitiallize: begin
				WE = 1;				// Write in random data
				on = 1;				// Start LFSR
				Address = count0;
				dataIn = data;
				if (count0 == 10'd164) begin
					nextState = halt;
					count0 = 0;
					count1 = 0;
				  Clear = 1;			// Clear the data of sum in hiddenlayer_top
				end
				else
				  count0++;
			end
			// For reading weight in test bench.
			readWeight: begin
				WE = 0;
				Clear = 0;
				inVal = in1[count0];
				if(dataOut) begin
      				weight = dataOut;
      				nextState = hiddenLayer;
  				end
  				else
  				  nextState = halt;
			end
			halt1: begin
				on = 0;
				out_hid = out0;
				Address = count0 + 8'd150 + count1*8'd5;
				nextState = readWeight1;
			end
			// The states above used to initiallize the weight.
			// ****************************************************************//
			// Hidden Layer for sum calculation
			hiddenLayer: begin // Calculate the output value of hiddenLayer
				AF_in = sum;
				out0[count1] = AF;
				if (count1 == 4) begin
				  nextState = halt1;
				  Clear = 1;
				  count0 = 0;
				  count1 = 0;
				end
				else begin
				  if (count0 == 29) begin
				    count1++;
				    count0 = 0;
				    Clear = 1;
				    nextState = halt;
				  end
				  else begin
				    count0++;
				    nextState = halt;
				  end
				end
			end
			outputLayer: begin
				AF_in = sum;
				out1[count1] = AF;
				if(count1 ==2) begin
					nextState = halt2;
				end
				else begin
					if(count0 == 4) begin
						count1++;
						count0 = 0;
						Clear = 1;
						nextState = halt1;
					end
					else begin
						count0++;
						nextState = halt1;
					end
				end
			end
			readWeight1: begin
				WE = 0;
				Clear = 0;
				inVal1 = out_hid[count0];
				if(dataOut) begin
      				weight = dataOut;
      				nextState = outputLayer;
  				end
				else
				  nextState = halt1;
			end
			halt2: begin
				Clear = 1;
				count0 = 0;
				count1 = 0;
				out_ann = out1;
				if(training)
					nextState = weightOptimize;
				else
					nextState = halt;
			end
			weightOptimize: begin //read weight first.
				WE = 0;
				Address = count0 + 8'd150 + count1*8'd5;
				if(dataOut) 
      				nextState = weightUpdate;
  				else
  				  nextState = weightOptimize;
			end
			weightUpdate: begin
				if(sign1[count1])
					dataIn = dataOut-delta1[count1];
				else
					dataIn = dataOut+delta1[count1];
				if(dataIn) 
      				nextState = writeWeight;
  				else if(dataIn == 0)
  				  nextState = writeWeight;
				else 
				  nextState = weightUpdate;
			end
			writeWeight: begin
			  WE = 1;
				if(count1 == 2) begin
					nextState = halt;
				end
				else begin
					if(count0 == 4)begin
						count1++;
						count0 = 0;
						nextState = weightOptimize;
					end
					else begin
						count0++;
						nextState = weightOptimize;
					end
				end
			end
		endcase
	end
	
	// The following sections are for output layer.
	// ******************************************************************
	// Get the error between calculated output and actual output.
	Subtraction sub1_0(out_ann_real[0],out_ann[0],out1_err[0],sign1[0]);
	Subtraction sub1_1(out_ann_real[1],out_ann[1],out1_err[1],sign1[1]);
	Subtraction sub1_2(out_ann_real[2],out_ann[2],out1_err[2],sign1[2]);
	
	SigmoidPrime sig1_0(out_ann[0],sig_prime_1[0]);
	SigmoidPrime sig1_1(out_ann[1],sig_prime_1[1]);
	SigmoidPrime sig1_2(out_ann[2],sig_prime_1[2]);
	
	// Calculate the value that need to change for weight1
	Delta delta1_0(out1_err[0],sig_prime_1[0],delta1[0]);
	Delta delta1_1(out1_err[1],sig_prime_1[1],delta1[1]);
	Delta delta1_2(out1_err[2],sig_prime_1[2],delta1[2]);
	
	// For hidden layer calculation.
	HiddenLayer_top getMul(Clock, Clear, weight, inVal, sum);
	ActivationFunc actFun(AF_in, AF);
	
	// For weight initiallize.
	LFSR rndnm(Clock, Rst, on, data);
	WeightRAM ram(Clock, Rst, dataIn, Address, WE, dataOut);
	
	
endmodule 