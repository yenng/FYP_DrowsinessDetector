module HiddenLayer(
	input Clock, WE,In,
	input [9:0] inVal[9:0],
	input [9:0] weight[9:0],
	output [1:0]outVal
);

integer i;
always@(posedge Clock)begin
end

endmodule
