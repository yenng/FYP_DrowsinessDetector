library verilog;
use verilog.vl_types.all;
entity Delta_tb is
end Delta_tb;
