library verilog;
use verilog.vl_types.all;
entity WeightInitiallize_tb is
end WeightInitiallize_tb;
