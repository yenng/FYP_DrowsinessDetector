library verilog;
use verilog.vl_types.all;
entity LFSR_tb is
end LFSR_tb;
