library verilog;
use verilog.vl_types.all;
entity WeighInitiallize_tb is
end WeighInitiallize_tb;
