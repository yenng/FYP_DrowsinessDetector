module DrowsinessDetector(
	input Clock,Rst,Start,
	input [9:0]in[0:9],
	output reg signed[9:0] weight,dataIn,
	output reg [9:0] outVal);
	
	//reg [639:0]testVal[0:479];
	
	// Slow Clock.
	reg Clock_slow;
	
	// For counter.
	reg [9:0]count0;		// The number that count in counter.
	reg [9:0]count1;
	reg startCounter0;		// To start the counter.
	reg startCounter1;
	wire stopCounter0;		// To stop the counter.
	wire stopCounter1;
	reg [9:0]max;			// Max value for counter.
	
	// For RAM to write/read weight. 
	reg WE;
	
	// The random data that generated by LFSR.
	reg signed[9:0] data;
	reg on;
	
	// The address of RAM to call the weight.
	reg [6:0] Address;
	
	// The variable that represent the state and nextState.
	reg [3:0] state;
	reg [3:0] nextState;
	
	// Parameter for the state.
	parameter 	halt = 0, weightInitiallize = 1, readWeight = 2, halt1 = 3, hiddenLayer_sum = 4,
	           hiddenLayer_AF = 5;
	
	// The variable for hidden layer.
	reg Clear;
	reg signed[9:0]sum;
	//reg [9:0]
	reg unsigned[9:0]inVal;
	
	always@(posedge Clock, negedge Rst) begin
		if(~Rst) begin
			state <= halt;
		end
		else begin
			state <= nextState;
		end
	end
	
	always@(stopCounter0, Start, state,data,sum) begin
		case(state)
		  // The following state is for weightInitiallize module.
			halt: begin
				startCounter0 = 0;	// Off and clear counter
				startCounter1 = 0;	// Off and clear counter
				on = 0;				// Off LFSR
				Clear = 1;
				if(Start)
					nextState = hiddenLayer_sum;
				else
					nextState = weightInitiallize;
			end
			weightInitiallize: begin
				WE = 1;				// Start counter
				on = 1;				// Start LFSR
				dataIn = data;
				max = 10'd65;
				startCounter0 = 1;
				if (stopCounter0) begin
					nextState = halt;
				end
			end
			// For reading weight in test bench.
			readWeight: begin
				WE = 0;
				on = 1;
				startCounter0 = 1;	// Start counter
			end
			halt1: begin
				startCounter0 = 0;	// Off and clear counter
				on = 0;
				Clear = 1;
				//nextState = readWeight;
			end
			// The states above used to initiallize the weight.
			// ****************************************************************//
			// Hidden Layer for sum calculation
			hiddenLayer_sum: begin // Calculate the sum of weight*in
				max = $size(in);
				startCounter0 = 1;
				startCounter1 = 1;
				Clear = 0;
				WE = 0;
				inVal = in[count0];
				Address = count0 + count1* 6'd10;
				outVal = sum;
				AF_in = sum;
				//weight = dataRead;
				if (stopCounter0) begin
					nextState = hiddenLayer_AF;
				end
			end
			// Hidden Layer for Activation Function.
			hiddenLayer_AF: begin
				Clear = 1;
				startCounter0 = 0;
				on = 0;
				outVal = AF;
				nextState = halt1;
			end
		endcase
	end
	
	// For a slower clock.
	clk_div createSlowClk(Clock, Clock_slow);
	
	// For hidden layer calculation.
	HiddenLayer_top getMul(Clock, Clear, weight, inVal, sum);
	ActivationFunc actFun(AF_in, AF);
	
	// For weight initiallize.
	LFSR rndnm(Clock, Rst, on, data);
	counter counter0(Clock, startCounter0, max, stopCounter0, count0);
	counter counter1(Clock_slow, startCounter1, 10'd10, stopCounter1, count1);
	WeightRAM ram(Clock, Rst, dataIn, Address, WE, weight);
	
	
endmodule 