library verilog;
use verilog.vl_types.all;
entity ActivationFunc_tb is
end ActivationFunc_tb;
